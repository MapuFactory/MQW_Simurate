* 40;Circuit4.ckt

.CIRCUITNAME "Circuit4"
.rootnamemap 40;Circuit4
.namemap
Z3=40;Circuit4;45
Z1=40;Circuit4;41
Z2=40;Circuit4;44
C6=40;Circuit4;100
Z4=40;Circuit4;46
C1=40;Circuit4;72
C2=40;Circuit4;74
L2=40;Circuit4;73
C4=40;Circuit4;88
L3=40;Circuit4;89
L4=40;Circuit4;90
C3=40;Circuit4;87
L6=40;Circuit4;99
L1=40;Circuit4;71
C5=40;Circuit4;112
L5=40;Circuit4;111
.endnamemap
.stringparam syslib = "C:\Program Files (x86)\Ansoft\DesignerSV2\syslib"
.stringparam userlib = "C:\Program Files (x86)\Ansoft\DesignerSV2\userlib"
.stringparam personallib = "C:\Users\kamei-lab\Documents\Ansoft\PersonalLib"
.stringparam projectdir = "C:\Users\kamei-lab\Desktop\miyata\text-20181004T040059Z-001\text\fig\designer"

*begin toplevel circuit
.param g1=0.629100000000000
.param g3=0.629100000000000
.param g2=0.970200000000000
.param g0=1
.param g4=1
.param Z0=50
.param w0={2*pi*1000000000.}
.param w1={2*pi*900000000}
.param w2={2*pi*1200000000.}
.param w3={2*pi*2300000000.}
.param w4={2*pi*2500000000.}
.param A1={w4 - w3 + w2 - w1}
.param B1={w1*w2*w3*w4/(w1*w2*w4 - w1*w2*w3 + w2*w3*w4 - w1*w3*w4)}
.param A2={(w2 - w3)*(w4 - w3)*(w2 + w4)*(w1 + w3)*(w1 - w2)*(w4 - w1)/(w1*w2*w4 - w1*w2*w3 + w2*w3*w4 - w1*w3*w4)/A1/A1}
.param B2={(w1*w2*w4 - w1*w2*w3 + w2*w3*w4 - w1*w3*w4)^2*A1/(w2 - w3)/(w4 - w3)/(w2 + w4)/(w1 + w3)/(w1 - w2)/(w4 - w1)}
.param J1=0.0100000000000000
.param J2=0.0100000000000000
.param J3=0.0100000000000000
.param J4={J1*J3/J2}
JINV:45 net_383 net_384 JINV={J3}
JINV:41 Port1 net_382 JINV={J1}
JINV:44 net_382 net_383 JINV={J2}
CAP:100 0 net_359 C={g3*Z0/B2*J1*J1*J3*J3/J2/J2} 
JINV:46 net_384 Port2 JINV={J4}
CAP:72 0 net_382 C={g1*Z0/A1*J1*J1} 
CAP:74 0 net_287 C={g1*Z0/B2*J1*J1} 
IND:73 net_287 net_382 L={1/g1/Z0/A2/J1/J1} 
CAP:88 0 net_304 C={g2/Z0/B2*J2*J2/J1/J1} 
IND:89 0 net_383 L={Z0/g2/B1*J1*J1/J2/J2} 
IND:90 net_304 net_383 L={Z0/g2/A2*J1*J1/J2/J2} 
CAP:87 0 net_383 C={g2/Z0/A1*J2*J2/J1/J1} 
IND:99 net_359 net_384 L={1/g3/Z0/A2/J1/J1/J3/J3*J2*J2} 
IND:71 0 net_382 L={1/g1/Z0/B1/J1/J1} 
CAP:112 0 net_384 C={g3*Z0/A1*J1*J1*J3*J3/J2/J2} 
IND:111 0 net_384 L={1/g3/Z0/B1/J1/J1/J3/J3*J2*J2} 
PORT:Port1 Port1 0 PNUM=1 rz={g0*Z0} iz=0Ohm 
PORT:Port2 Port2 0 PNUM=2 rz={g4*Z0} iz=0Ohm 


*end toplevel circuit
.nwa:"NWA1"
+ F=LIN 1MHz 10GHz 1MHz
+ SWPORD = {F}
+ SolutionFile="C:\Users\kamei-lab\Documents\Ansoft\temp\Project1.results\Circuit4_NWA1_61_U4_Circuit4_401_398\Circuit4_NWA1_61_U4_Circuit4_401_398.sol"

.end
